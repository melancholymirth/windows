module inverter(input in, output out);

	assign in = ~out;

endmodule