/* This is our control unit.
It contains our state machine, which has 3 states:
1) HALT state
2) COUNT (for #0-6) --> implement the ADD operation (depending on 'M')
3) COUNT for #7 --> implement the ADD/SUBTRACT operation (depending on 'M')
*/
module control();

endmodule
