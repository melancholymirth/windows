module multiplier_8bit(
		
		input logic enable, clk, reset,
		output logic [7:0] out);
		
		
		counter myCounter(.*);
		
		
endmodule